package shared_pkg;
int unsigned error_count;
int unsigned correct_count;
bit test_done;
endpackage
 